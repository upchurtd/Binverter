library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


ENTITY VGA IS
PORT(
	CLOCK_24: IN STD_LOGIC_VECTOR(1 downto 0);
	VGA_HS,VGA_VS:OUT STD_LOGIC;
	--SW: STD_LOGIC_VECTOR(1 downto 0);
	--KEY: STD_LOGIC_VECTOR(3 DOWNTO 0);
	VGA_R,VGA_B,VGA_G: OUT STD_LOGIC_VECTOR(3 downto 0)
);
END VGA;


ARCHITECTURE MAIN OF VGA IS
	--SIGNAL VGACLK,RESET:STD_LOGIC;

COMPONENT SYNC IS
 PORT(
	CLK: IN STD_LOGIC;
	HSYNC: OUT STD_LOGIC;
	VSYNC: OUT STD_LOGIC;
	R, G, B: OUT STD_LOGIC_VECTOR(3 downto 0);
	--KEYS: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
   --S: IN STD_LOGIC_VECTOR(1 downto 0)
	);
END COMPONENT SYNC;



    component pll is
        port (
            clkout_clk : out std_logic;        -- clk
            clkin_clk  : in  std_logic := 'X'; -- clk
            rst_reset  : in  std_logic := 'X'  -- reset
        );
	 END COMPONENT pll;
 BEGIN
 
 --C: pll PORT MAP (VGACLK,CLOCK_24(0),RESET);
 --C1: SYNC PORT MAP(VGACLK,VGA_HS,VGA_VS,VGA_R,VGA_G,VGA_B,KEY,SW);
 C1: SYNC PORT MAP(VGACLK,VGA_HS,VGA_VS,VGA_R,VGA_G,VGA_B);
 
 END MAIN;